module top_module(
	input a,b,c,d,e,
	output [24:0] out
);
	wire [24:0] t1,t2;
	assign t1 = {{5{a}},{5{b}},{5{c}},{5{d}},{5{e}}};
	assign t2 = {5{a,b,c,d,e}};
	assign out = ~ t1 ^ t2;

endmodule
